// mySystem.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module mySystem (
		input  wire        alt_vip_cl_cvo_0_clocked_video_vid_clk,                      //                  alt_vip_cl_cvo_0_clocked_video.vid_clk
		output wire [23:0] alt_vip_cl_cvo_0_clocked_video_vid_data,                     //                                                .vid_data
		output wire        alt_vip_cl_cvo_0_clocked_video_underflow,                    //                                                .underflow
		output wire        alt_vip_cl_cvo_0_clocked_video_vid_datavalid,                //                                                .vid_datavalid
		output wire        alt_vip_cl_cvo_0_clocked_video_vid_v_sync,                   //                                                .vid_v_sync
		output wire        alt_vip_cl_cvo_0_clocked_video_vid_h_sync,                   //                                                .vid_h_sync
		output wire        alt_vip_cl_cvo_0_clocked_video_vid_f,                        //                                                .vid_f
		output wire        alt_vip_cl_cvo_0_clocked_video_vid_h,                        //                                                .vid_h
		output wire        alt_vip_cl_cvo_0_clocked_video_vid_v,                        //                                                .vid_v
		input  wire        alt_vip_cti_0_clocked_video_vid_clk,                         //                     alt_vip_cti_0_clocked_video.vid_clk
		input  wire [23:0] alt_vip_cti_0_clocked_video_vid_data,                        //                                                .vid_data
		output wire        alt_vip_cti_0_clocked_video_overflow,                        //                                                .overflow
		input  wire        alt_vip_cti_0_clocked_video_vid_datavalid,                   //                                                .vid_datavalid
		input  wire        alt_vip_cti_0_clocked_video_vid_locked,                      //                                                .vid_locked
		input  wire        alt_vip_cti_0_clocked_video_vid_v_sync,                      //                                                .vid_v_sync
		input  wire        alt_vip_cti_0_clocked_video_vid_h_sync,                      //                                                .vid_h_sync
		input  wire        alt_vip_cti_0_clocked_video_vid_f,                           //                                                .vid_f
		input  wire        clk_clk,                                                     //                                             clk.clk
		output wire [1:0]  pio_0_external_connection_export,                            //                       pio_0_external_connection.export
		input  wire        reset_reset_n,                                               //                                           reset.reset_n
		input  wire        uart_0_external_connection_rxd,                              //                      uart_0_external_connection.rxd
		output wire        uart_0_external_connection_txd,                              //                                                .txd
		output wire [12:0] w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if_sdram_addr,  // w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if.sdram_addr
		output wire [1:0]  w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if_sdram_ba,    //                                                .sdram_ba
		output wire        w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if_sdram_cas_n, //                                                .sdram_cas_n
		output wire        w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if_sdram_cke,   //                                                .sdram_cke
		output wire        w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if_sdram_cs_n,  //                                                .sdram_cs_n
		inout  wire [15:0] w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if_sdram_dq,    //                                                .sdram_dq
		output wire [1:0]  w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if_sdram_dqm,   //                                                .sdram_dqm
		output wire        w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if_sdram_ras_n, //                                                .sdram_ras_n
		output wire        w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if_sdram_we_n   //                                                .sdram_we_n
	);

	wire         alt_vip_cl_mixer_0_dout_valid;                                                         // alt_vip_cl_mixer_0:dout_valid -> alt_vip_cl_cvo_0:din_valid
	wire  [23:0] alt_vip_cl_mixer_0_dout_data;                                                          // alt_vip_cl_mixer_0:dout_data -> alt_vip_cl_cvo_0:din_data
	wire         alt_vip_cl_mixer_0_dout_ready;                                                         // alt_vip_cl_cvo_0:din_ready -> alt_vip_cl_mixer_0:dout_ready
	wire         alt_vip_cl_mixer_0_dout_startofpacket;                                                 // alt_vip_cl_mixer_0:dout_startofpacket -> alt_vip_cl_cvo_0:din_startofpacket
	wire         alt_vip_cl_mixer_0_dout_endofpacket;                                                   // alt_vip_cl_mixer_0:dout_endofpacket -> alt_vip_cl_cvo_0:din_endofpacket
	wire         alt_vip_cl_tpg_0_dout_valid;                                                           // alt_vip_cl_tpg_0:dout_valid -> main_scaler:din_valid
	wire  [23:0] alt_vip_cl_tpg_0_dout_data;                                                            // alt_vip_cl_tpg_0:dout_data -> main_scaler:din_data
	wire         alt_vip_cl_tpg_0_dout_ready;                                                           // main_scaler:din_ready -> alt_vip_cl_tpg_0:dout_ready
	wire         alt_vip_cl_tpg_0_dout_startofpacket;                                                   // alt_vip_cl_tpg_0:dout_startofpacket -> main_scaler:din_startofpacket
	wire         alt_vip_cl_tpg_0_dout_endofpacket;                                                     // alt_vip_cl_tpg_0:dout_endofpacket -> main_scaler:din_endofpacket
	wire         main_scaler_dout_valid;                                                                // main_scaler:dout_valid -> alt_vip_cl_vfb_0:din_valid
	wire  [23:0] main_scaler_dout_data;                                                                 // main_scaler:dout_data -> alt_vip_cl_vfb_0:din_data
	wire         main_scaler_dout_ready;                                                                // alt_vip_cl_vfb_0:din_ready -> main_scaler:dout_ready
	wire         main_scaler_dout_startofpacket;                                                        // main_scaler:dout_startofpacket -> alt_vip_cl_vfb_0:din_startofpacket
	wire         main_scaler_dout_endofpacket;                                                          // main_scaler:dout_endofpacket -> alt_vip_cl_vfb_0:din_endofpacket
	wire         alt_vip_cl_vfb_0_dout_valid;                                                           // alt_vip_cl_vfb_0:dout_valid -> alt_vip_cl_mixer_0:din0_valid
	wire  [23:0] alt_vip_cl_vfb_0_dout_data;                                                            // alt_vip_cl_vfb_0:dout_data -> alt_vip_cl_mixer_0:din0_data
	wire         alt_vip_cl_vfb_0_dout_ready;                                                           // alt_vip_cl_mixer_0:din0_ready -> alt_vip_cl_vfb_0:dout_ready
	wire         alt_vip_cl_vfb_0_dout_startofpacket;                                                   // alt_vip_cl_vfb_0:dout_startofpacket -> alt_vip_cl_mixer_0:din0_startofpacket
	wire         alt_vip_cl_vfb_0_dout_endofpacket;                                                     // alt_vip_cl_vfb_0:dout_endofpacket -> alt_vip_cl_mixer_0:din0_endofpacket
	wire         alt_vip_cti_0_dout_valid;                                                              // alt_vip_cti_0:is_valid -> alt_vip_cl_mixer_0:din1_valid
	wire  [23:0] alt_vip_cti_0_dout_data;                                                               // alt_vip_cti_0:is_data -> alt_vip_cl_mixer_0:din1_data
	wire         alt_vip_cti_0_dout_ready;                                                              // alt_vip_cl_mixer_0:din1_ready -> alt_vip_cti_0:is_ready
	wire         alt_vip_cti_0_dout_startofpacket;                                                      // alt_vip_cti_0:is_sop -> alt_vip_cl_mixer_0:din1_startofpacket
	wire         alt_vip_cti_0_dout_endofpacket;                                                        // alt_vip_cti_0:is_eop -> alt_vip_cl_mixer_0:din1_endofpacket
	wire  [31:0] nios2_gen2_0_data_master_readdata;                                                     // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                                                  // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                                                  // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [14:0] nios2_gen2_0_data_master_address;                                                      // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                                                   // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                                         // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                                                        // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                                                    // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                                              // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                                           // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [14:0] nios2_gen2_0_instruction_master_address;                                               // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                                                  // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire  [31:0] mm_interconnect_0_alt_vip_cl_mixer_0_control_readdata;                                 // alt_vip_cl_mixer_0:control_readdata -> mm_interconnect_0:alt_vip_cl_mixer_0_control_readdata
	wire         mm_interconnect_0_alt_vip_cl_mixer_0_control_waitrequest;                              // alt_vip_cl_mixer_0:control_waitrequest -> mm_interconnect_0:alt_vip_cl_mixer_0_control_waitrequest
	wire   [6:0] mm_interconnect_0_alt_vip_cl_mixer_0_control_address;                                  // mm_interconnect_0:alt_vip_cl_mixer_0_control_address -> alt_vip_cl_mixer_0:control_address
	wire         mm_interconnect_0_alt_vip_cl_mixer_0_control_read;                                     // mm_interconnect_0:alt_vip_cl_mixer_0_control_read -> alt_vip_cl_mixer_0:control_read
	wire   [3:0] mm_interconnect_0_alt_vip_cl_mixer_0_control_byteenable;                               // mm_interconnect_0:alt_vip_cl_mixer_0_control_byteenable -> alt_vip_cl_mixer_0:control_byteenable
	wire         mm_interconnect_0_alt_vip_cl_mixer_0_control_readdatavalid;                            // alt_vip_cl_mixer_0:control_readdatavalid -> mm_interconnect_0:alt_vip_cl_mixer_0_control_readdatavalid
	wire         mm_interconnect_0_alt_vip_cl_mixer_0_control_write;                                    // mm_interconnect_0:alt_vip_cl_mixer_0_control_write -> alt_vip_cl_mixer_0:control_write
	wire  [31:0] mm_interconnect_0_alt_vip_cl_mixer_0_control_writedata;                                // mm_interconnect_0:alt_vip_cl_mixer_0_control_writedata -> alt_vip_cl_mixer_0:control_writedata
	wire  [31:0] mm_interconnect_0_main_scaler_control_readdata;                                        // main_scaler:control_readdata -> mm_interconnect_0:main_scaler_control_readdata
	wire         mm_interconnect_0_main_scaler_control_waitrequest;                                     // main_scaler:control_waitrequest -> mm_interconnect_0:main_scaler_control_waitrequest
	wire   [6:0] mm_interconnect_0_main_scaler_control_address;                                         // mm_interconnect_0:main_scaler_control_address -> main_scaler:control_address
	wire         mm_interconnect_0_main_scaler_control_read;                                            // mm_interconnect_0:main_scaler_control_read -> main_scaler:control_read
	wire   [3:0] mm_interconnect_0_main_scaler_control_byteenable;                                      // mm_interconnect_0:main_scaler_control_byteenable -> main_scaler:control_byteenable
	wire         mm_interconnect_0_main_scaler_control_readdatavalid;                                   // main_scaler:control_readdatavalid -> mm_interconnect_0:main_scaler_control_readdatavalid
	wire         mm_interconnect_0_main_scaler_control_write;                                           // mm_interconnect_0:main_scaler_control_write -> main_scaler:control_write
	wire  [31:0] mm_interconnect_0_main_scaler_control_writedata;                                       // mm_interconnect_0:main_scaler_control_writedata -> main_scaler:control_writedata
	wire  [15:0] mm_interconnect_0_alt_vip_cti_0_control_readdata;                                      // alt_vip_cti_0:av_readdata -> mm_interconnect_0:alt_vip_cti_0_control_readdata
	wire   [3:0] mm_interconnect_0_alt_vip_cti_0_control_address;                                       // mm_interconnect_0:alt_vip_cti_0_control_address -> alt_vip_cti_0:av_address
	wire         mm_interconnect_0_alt_vip_cti_0_control_read;                                          // mm_interconnect_0:alt_vip_cti_0_control_read -> alt_vip_cti_0:av_read
	wire         mm_interconnect_0_alt_vip_cti_0_control_write;                                         // mm_interconnect_0:alt_vip_cti_0_control_write -> alt_vip_cti_0:av_write
	wire  [15:0] mm_interconnect_0_alt_vip_cti_0_control_writedata;                                     // mm_interconnect_0:alt_vip_cti_0_control_writedata -> alt_vip_cti_0:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;                               // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;                            // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;                            // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;                                // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;                                   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;                             // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;                                  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;                              // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                                      // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                                        // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [10:0] mm_interconnect_0_onchip_memory2_0_s1_address;                                         // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                                      // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                                           // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                                       // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                                           // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_pio_0_s1_chipselect;                                                 // mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;                                                   // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;                                                    // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_pio_0_s1_write;                                                      // mm_interconnect_0:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;                                                  // mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	wire         mm_interconnect_0_uart_0_s1_chipselect;                                                // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;                                                  // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;                                                   // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_read;                                                      // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire         mm_interconnect_0_uart_0_s1_begintransfer;                                             // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_uart_0_s1_write;                                                     // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;                                                 // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire         alt_vip_cl_vfb_0_mem_master_rd_waitrequest;                                            // mm_interconnect_1:alt_vip_cl_vfb_0_mem_master_rd_waitrequest -> alt_vip_cl_vfb_0:mem_master_rd_waitrequest
	wire  [31:0] alt_vip_cl_vfb_0_mem_master_rd_readdata;                                               // mm_interconnect_1:alt_vip_cl_vfb_0_mem_master_rd_readdata -> alt_vip_cl_vfb_0:mem_master_rd_readdata
	wire  [31:0] alt_vip_cl_vfb_0_mem_master_rd_address;                                                // alt_vip_cl_vfb_0:mem_master_rd_address -> mm_interconnect_1:alt_vip_cl_vfb_0_mem_master_rd_address
	wire         alt_vip_cl_vfb_0_mem_master_rd_read;                                                   // alt_vip_cl_vfb_0:mem_master_rd_read -> mm_interconnect_1:alt_vip_cl_vfb_0_mem_master_rd_read
	wire         alt_vip_cl_vfb_0_mem_master_rd_readdatavalid;                                          // mm_interconnect_1:alt_vip_cl_vfb_0_mem_master_rd_readdatavalid -> alt_vip_cl_vfb_0:mem_master_rd_readdatavalid
	wire   [5:0] alt_vip_cl_vfb_0_mem_master_rd_burstcount;                                             // alt_vip_cl_vfb_0:mem_master_rd_burstcount -> mm_interconnect_1:alt_vip_cl_vfb_0_mem_master_rd_burstcount
	wire         alt_vip_cl_vfb_0_mem_master_wr_waitrequest;                                            // mm_interconnect_1:alt_vip_cl_vfb_0_mem_master_wr_waitrequest -> alt_vip_cl_vfb_0:mem_master_wr_waitrequest
	wire  [31:0] alt_vip_cl_vfb_0_mem_master_wr_address;                                                // alt_vip_cl_vfb_0:mem_master_wr_address -> mm_interconnect_1:alt_vip_cl_vfb_0_mem_master_wr_address
	wire   [3:0] alt_vip_cl_vfb_0_mem_master_wr_byteenable;                                             // alt_vip_cl_vfb_0:mem_master_wr_byteenable -> mm_interconnect_1:alt_vip_cl_vfb_0_mem_master_wr_byteenable
	wire         alt_vip_cl_vfb_0_mem_master_wr_write;                                                  // alt_vip_cl_vfb_0:mem_master_wr_write -> mm_interconnect_1:alt_vip_cl_vfb_0_mem_master_wr_write
	wire  [31:0] alt_vip_cl_vfb_0_mem_master_wr_writedata;                                              // alt_vip_cl_vfb_0:mem_master_wr_writedata -> mm_interconnect_1:alt_vip_cl_vfb_0_mem_master_wr_writedata
	wire   [5:0] alt_vip_cl_vfb_0_mem_master_wr_burstcount;                                             // alt_vip_cl_vfb_0:mem_master_wr_burstcount -> mm_interconnect_1:alt_vip_cl_vfb_0_mem_master_wr_burstcount
	wire         mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_chipselect;    // mm_interconnect_1:W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0_chipselect -> W9825G6KH_SDRAMController_125MHz_CL3_0:az_cs
	wire  [15:0] mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_readdata;      // W9825G6KH_SDRAMController_125MHz_CL3_0:za_data -> mm_interconnect_1:W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0_readdata
	wire         mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_waitrequest;   // W9825G6KH_SDRAMController_125MHz_CL3_0:za_waitrequest -> mm_interconnect_1:W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0_waitrequest
	wire  [23:0] mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_address;       // mm_interconnect_1:W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0_address -> W9825G6KH_SDRAMController_125MHz_CL3_0:az_addr
	wire         mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_read;          // mm_interconnect_1:W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0_read -> W9825G6KH_SDRAMController_125MHz_CL3_0:az_rd_n
	wire   [1:0] mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_byteenable;    // mm_interconnect_1:W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0_byteenable -> W9825G6KH_SDRAMController_125MHz_CL3_0:az_be_n
	wire         mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_readdatavalid; // W9825G6KH_SDRAMController_125MHz_CL3_0:za_valid -> mm_interconnect_1:W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0_readdatavalid
	wire         mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_write;         // mm_interconnect_1:W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0_write -> W9825G6KH_SDRAMController_125MHz_CL3_0:az_wr_n
	wire  [15:0] mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_writedata;     // mm_interconnect_1:W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0_writedata -> W9825G6KH_SDRAMController_125MHz_CL3_0:az_data
	wire         irq_mapper_receiver0_irq;                                                              // uart_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                              // alt_vip_cti_0:status_update_int -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                                                  // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                                                        // rst_controller:reset_out -> [W9825G6KH_SDRAMController_125MHz_CL3_0:reset_n, alt_vip_cl_cvo_0:main_reset_reset, alt_vip_cl_mixer_0:main_reset_reset, alt_vip_cl_tpg_0:main_reset, alt_vip_cl_vfb_0:main_reset, alt_vip_cl_vfb_0:mem_reset, alt_vip_cti_0:rst, irq_mapper:reset, main_scaler:main_reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:alt_vip_cl_vfb_0_mem_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, pio_0:reset_n, rst_translator:in_reset, uart_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                                                    // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	W9825G6KH_SDRAMController_125MHz_CL3 w9825g6kh_sdramcontroller_125mhz_cl3_0 (
		.az_addr        (mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_address),       // avalon_slave_0.address
		.az_be_n        (~mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_byteenable),   //               .byteenable_n
		.az_cs          (mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_chipselect),    //               .chipselect
		.az_data        (mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_writedata),     //               .writedata
		.az_rd_n        (~mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_read),         //               .read_n
		.az_wr_n        (~mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_write),        //               .write_n
		.za_data        (mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_readdata),      //               .readdata
		.za_valid       (mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_readdatavalid), //               .readdatavalid
		.za_waitrequest (mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_waitrequest),   //               .waitrequest
		.clk            (clk_clk),                                                                               //          clock.clk
		.reset_n        (~rst_controller_reset_out_reset),                                                       //          reset.reset_n
		.zs_addr        (w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if_sdram_addr),                            //       sdram_if.sdram_addr
		.zs_ba          (w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if_sdram_ba),                              //               .sdram_ba
		.zs_cas_n       (w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if_sdram_cas_n),                           //               .sdram_cas_n
		.zs_cke         (w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if_sdram_cke),                             //               .sdram_cke
		.zs_cs_n        (w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if_sdram_cs_n),                            //               .sdram_cs_n
		.zs_dq          (w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if_sdram_dq),                              //               .sdram_dq
		.zs_dqm         (w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if_sdram_dqm),                             //               .sdram_dqm
		.zs_ras_n       (w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if_sdram_ras_n),                           //               .sdram_ras_n
		.zs_we_n        (w9825g6kh_sdramcontroller_125mhz_cl3_0_sdram_if_sdram_we_n)                             //               .sdram_we_n
	);

	mySystem_alt_vip_cl_cvo_0 #(
		.BPS                           (8),
		.NUMBER_OF_COLOUR_PLANES       (3),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (640),
		.V_ACTIVE_LINES                (480),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (640),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (639),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.ACCEPT_SYNC                   (0),
		.COUNT_STEP_IS_PIP_VALUE       (0),
		.LOW_LATENCY                   (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (96),
		.H_FRONT_PORCH                 (16),
		.H_BACK_PORCH                  (48),
		.V_SYNC_LENGTH                 (2),
		.V_FRONT_PORCH                 (11),
		.V_BACK_PORCH                  (31),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0),
		.PIXELS_IN_PARALLEL            (1),
		.SRC_WIDTH                     (8),
		.DST_WIDTH                     (8),
		.CONTEXT_WIDTH                 (8),
		.TASK_WIDTH                    (8)
	) alt_vip_cl_cvo_0 (
		.clocked_video_vid_clk       (alt_vip_cl_cvo_0_clocked_video_vid_clk),       // clocked_video.vid_clk
		.clocked_video_vid_data      (alt_vip_cl_cvo_0_clocked_video_vid_data),      //              .vid_data
		.clocked_video_underflow     (alt_vip_cl_cvo_0_clocked_video_underflow),     //              .underflow
		.clocked_video_vid_datavalid (alt_vip_cl_cvo_0_clocked_video_vid_datavalid), //              .vid_datavalid
		.clocked_video_vid_v_sync    (alt_vip_cl_cvo_0_clocked_video_vid_v_sync),    //              .vid_v_sync
		.clocked_video_vid_h_sync    (alt_vip_cl_cvo_0_clocked_video_vid_h_sync),    //              .vid_h_sync
		.clocked_video_vid_f         (alt_vip_cl_cvo_0_clocked_video_vid_f),         //              .vid_f
		.clocked_video_vid_h         (alt_vip_cl_cvo_0_clocked_video_vid_h),         //              .vid_h
		.clocked_video_vid_v         (alt_vip_cl_cvo_0_clocked_video_vid_v),         //              .vid_v
		.main_clock_clk              (clk_clk),                                      //    main_clock.clk
		.main_reset_reset            (rst_controller_reset_out_reset),               //    main_reset.reset
		.din_data                    (alt_vip_cl_mixer_0_dout_data),                 //           din.data
		.din_valid                   (alt_vip_cl_mixer_0_dout_valid),                //              .valid
		.din_startofpacket           (alt_vip_cl_mixer_0_dout_startofpacket),        //              .startofpacket
		.din_endofpacket             (alt_vip_cl_mixer_0_dout_endofpacket),          //              .endofpacket
		.din_ready                   (alt_vip_cl_mixer_0_dout_ready)                 //              .ready
	);

	mySystem_alt_vip_cl_mixer_0 #(
		.BITS_PER_SYMBOL              (8),
		.NUMBER_OF_COLOR_PLANES       (2),
		.COLOR_PLANES_ARE_IN_PARALLEL (1),
		.PIXELS_IN_PARALLEL           (1),
		.MAX_WIDTH                    (640),
		.MAX_HEIGHT                   (480),
		.IS_422                       (1),
		.LIMITED_READBACK             (0),
		.LOW_LATENCY_MODE             (0),
		.DATA_PIPELINE_STAGES         (0),
		.USER_PACKET_SUPPORT          ("DISCARD"),
		.USER_PACKET_FIFO_DEPTH       (0)
	) alt_vip_cl_mixer_0 (
		.main_clock_clk        (clk_clk),                                                    // main_clock.clk
		.main_reset_reset      (rst_controller_reset_out_reset),                             // main_reset.reset
		.din0_data             (alt_vip_cl_vfb_0_dout_data),                                 //       din0.data
		.din0_valid            (alt_vip_cl_vfb_0_dout_valid),                                //           .valid
		.din0_startofpacket    (alt_vip_cl_vfb_0_dout_startofpacket),                        //           .startofpacket
		.din0_endofpacket      (alt_vip_cl_vfb_0_dout_endofpacket),                          //           .endofpacket
		.din0_ready            (alt_vip_cl_vfb_0_dout_ready),                                //           .ready
		.din1_data             (alt_vip_cti_0_dout_data),                                    //       din1.data
		.din1_valid            (alt_vip_cti_0_dout_valid),                                   //           .valid
		.din1_startofpacket    (alt_vip_cti_0_dout_startofpacket),                           //           .startofpacket
		.din1_endofpacket      (alt_vip_cti_0_dout_endofpacket),                             //           .endofpacket
		.din1_ready            (alt_vip_cti_0_dout_ready),                                   //           .ready
		.dout_data             (alt_vip_cl_mixer_0_dout_data),                               //       dout.data
		.dout_valid            (alt_vip_cl_mixer_0_dout_valid),                              //           .valid
		.dout_startofpacket    (alt_vip_cl_mixer_0_dout_startofpacket),                      //           .startofpacket
		.dout_endofpacket      (alt_vip_cl_mixer_0_dout_endofpacket),                        //           .endofpacket
		.dout_ready            (alt_vip_cl_mixer_0_dout_ready),                              //           .ready
		.control_address       (mm_interconnect_0_alt_vip_cl_mixer_0_control_address),       //    control.address
		.control_byteenable    (mm_interconnect_0_alt_vip_cl_mixer_0_control_byteenable),    //           .byteenable
		.control_write         (mm_interconnect_0_alt_vip_cl_mixer_0_control_write),         //           .write
		.control_writedata     (mm_interconnect_0_alt_vip_cl_mixer_0_control_writedata),     //           .writedata
		.control_read          (mm_interconnect_0_alt_vip_cl_mixer_0_control_read),          //           .read
		.control_readdata      (mm_interconnect_0_alt_vip_cl_mixer_0_control_readdata),      //           .readdata
		.control_readdatavalid (mm_interconnect_0_alt_vip_cl_mixer_0_control_readdatavalid), //           .readdatavalid
		.control_waitrequest   (mm_interconnect_0_alt_vip_cl_mixer_0_control_waitrequest)    //           .waitrequest
	);

	mySystem_alt_vip_cl_tpg_0 #(
		.PIXELS_IN_PARALLEL (1)
	) alt_vip_cl_tpg_0 (
		.main_clock         (clk_clk),                             // main_clock.clk
		.main_reset         (rst_controller_reset_out_reset),      // main_reset.reset
		.dout_data          (alt_vip_cl_tpg_0_dout_data),          //       dout.data
		.dout_valid         (alt_vip_cl_tpg_0_dout_valid),         //           .valid
		.dout_startofpacket (alt_vip_cl_tpg_0_dout_startofpacket), //           .startofpacket
		.dout_endofpacket   (alt_vip_cl_tpg_0_dout_endofpacket),   //           .endofpacket
		.dout_ready         (alt_vip_cl_tpg_0_dout_ready)          //           .ready
	);

	mySystem_alt_vip_cl_vfb_0 #(
		.BITS_PER_SYMBOL              (8),
		.NUMBER_OF_COLOR_PLANES       (3),
		.COLOR_PLANES_ARE_IN_PARALLEL (1),
		.PIXELS_IN_PARALLEL           (1),
		.READY_LATENCY                (1),
		.MAX_WIDTH                    (640),
		.MAX_HEIGHT                   (480),
		.CLOCKS_ARE_SEPARATE          (1),
		.MEM_PORT_WIDTH               (32),
		.MEM_BASE_ADDR                (0),
		.BURST_ALIGNMENT              (1),
		.WRITE_FIFO_DEPTH             (64),
		.WRITE_BURST_TARGET           (32),
		.READ_FIFO_DEPTH              (64),
		.READ_BURST_TARGET            (32),
		.WRITER_RUNTIME_CONTROL       (0),
		.READER_RUNTIME_CONTROL       (0),
		.IS_FRAME_WRITER              (0),
		.IS_FRAME_READER              (0),
		.DROP_FRAMES                  (0),
		.REPEAT_FRAMES                (0),
		.DROP_REPEAT_USER             (0),
		.INTERLACED_SUPPORT           (0),
		.CONTROLLED_DROP_REPEAT       (0),
		.DROP_INVALID_FIELDS          (0),
		.MULTI_FRAME_DELAY            (1),
		.IS_SYNC_MASTER               (0),
		.IS_SYNC_SLAVE                (0),
		.LINE_BASED_BUFFERING         (0),
		.PRIORITIZE_FMAX              (0),
		.USER_PACKETS_MAX_STORAGE     (0),
		.MAX_SYMBOLS_PER_PACKET       (10),
		.NUM_BUFFERS                  (2)
	) alt_vip_cl_vfb_0 (
		.main_clock                  (clk_clk),                                      //    main_clock.clk
		.main_reset                  (rst_controller_reset_out_reset),               //    main_reset.reset
		.mem_clock                   (clk_clk),                                      //     mem_clock.clk
		.mem_reset                   (rst_controller_reset_out_reset),               //     mem_reset.reset
		.din_data                    (main_scaler_dout_data),                        //           din.data
		.din_valid                   (main_scaler_dout_valid),                       //              .valid
		.din_startofpacket           (main_scaler_dout_startofpacket),               //              .startofpacket
		.din_endofpacket             (main_scaler_dout_endofpacket),                 //              .endofpacket
		.din_ready                   (main_scaler_dout_ready),                       //              .ready
		.mem_master_wr_address       (alt_vip_cl_vfb_0_mem_master_wr_address),       // mem_master_wr.address
		.mem_master_wr_burstcount    (alt_vip_cl_vfb_0_mem_master_wr_burstcount),    //              .burstcount
		.mem_master_wr_waitrequest   (alt_vip_cl_vfb_0_mem_master_wr_waitrequest),   //              .waitrequest
		.mem_master_wr_write         (alt_vip_cl_vfb_0_mem_master_wr_write),         //              .write
		.mem_master_wr_writedata     (alt_vip_cl_vfb_0_mem_master_wr_writedata),     //              .writedata
		.mem_master_wr_byteenable    (alt_vip_cl_vfb_0_mem_master_wr_byteenable),    //              .byteenable
		.dout_data                   (alt_vip_cl_vfb_0_dout_data),                   //          dout.data
		.dout_valid                  (alt_vip_cl_vfb_0_dout_valid),                  //              .valid
		.dout_startofpacket          (alt_vip_cl_vfb_0_dout_startofpacket),          //              .startofpacket
		.dout_endofpacket            (alt_vip_cl_vfb_0_dout_endofpacket),            //              .endofpacket
		.dout_ready                  (alt_vip_cl_vfb_0_dout_ready),                  //              .ready
		.mem_master_rd_address       (alt_vip_cl_vfb_0_mem_master_rd_address),       // mem_master_rd.address
		.mem_master_rd_burstcount    (alt_vip_cl_vfb_0_mem_master_rd_burstcount),    //              .burstcount
		.mem_master_rd_waitrequest   (alt_vip_cl_vfb_0_mem_master_rd_waitrequest),   //              .waitrequest
		.mem_master_rd_read          (alt_vip_cl_vfb_0_mem_master_rd_read),          //              .read
		.mem_master_rd_readdata      (alt_vip_cl_vfb_0_mem_master_rd_readdata),      //              .readdata
		.mem_master_rd_readdatavalid (alt_vip_cl_vfb_0_mem_master_rd_readdatavalid)  //              .readdatavalid
	);

	alt_vipcti131_Vid2IS #(
		.BPS                           (8),
		.NUMBER_OF_COLOUR_PLANES       (3),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.SYNC_TO                       (2),
		.USE_EMBEDDED_SYNCS            (0),
		.ADD_DATA_ENABLE_SIGNAL        (0),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.USE_STD                       (0),
		.STD_WIDTH                     (1),
		.GENERATE_ANC                  (0),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS_F0            (1920),
		.V_ACTIVE_LINES_F0             (1080),
		.V_ACTIVE_LINES_F1             (32),
		.FIFO_DEPTH                    (1920),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (1),
		.GENERATE_SYNC                 (0)
	) alt_vip_cti_0 (
		.is_clk            (clk_clk),                                           //        is_clk_rst.clk
		.rst               (rst_controller_reset_out_reset),                    //  is_clk_rst_reset.reset
		.av_address        (mm_interconnect_0_alt_vip_cti_0_control_address),   //           control.address
		.av_read           (mm_interconnect_0_alt_vip_cti_0_control_read),      //                  .read
		.av_readdata       (mm_interconnect_0_alt_vip_cti_0_control_readdata),  //                  .readdata
		.av_write          (mm_interconnect_0_alt_vip_cti_0_control_write),     //                  .write
		.av_writedata      (mm_interconnect_0_alt_vip_cti_0_control_writedata), //                  .writedata
		.status_update_int (irq_mapper_receiver1_irq),                          // status_update_irq.irq
		.is_data           (alt_vip_cti_0_dout_data),                           //              dout.data
		.is_valid          (alt_vip_cti_0_dout_valid),                          //                  .valid
		.is_ready          (alt_vip_cti_0_dout_ready),                          //                  .ready
		.is_sop            (alt_vip_cti_0_dout_startofpacket),                  //                  .startofpacket
		.is_eop            (alt_vip_cti_0_dout_endofpacket),                    //                  .endofpacket
		.vid_clk           (alt_vip_cti_0_clocked_video_vid_clk),               //     clocked_video.export
		.vid_data          (alt_vip_cti_0_clocked_video_vid_data),              //                  .export
		.overflow          (alt_vip_cti_0_clocked_video_overflow),              //                  .export
		.vid_datavalid     (alt_vip_cti_0_clocked_video_vid_datavalid),         //                  .export
		.vid_locked        (alt_vip_cti_0_clocked_video_vid_locked),            //                  .export
		.vid_v_sync        (alt_vip_cti_0_clocked_video_vid_v_sync),            //                  .export
		.vid_h_sync        (alt_vip_cti_0_clocked_video_vid_h_sync),            //                  .export
		.vid_f             (alt_vip_cti_0_clocked_video_vid_f)                  //                  .export
	);

	mySystem_main_scaler main_scaler (
		.main_clock            (clk_clk),                                             // main_clock.clk
		.main_reset            (rst_controller_reset_out_reset),                      // main_reset.reset
		.din_data              (alt_vip_cl_tpg_0_dout_data),                          //        din.data
		.din_valid             (alt_vip_cl_tpg_0_dout_valid),                         //           .valid
		.din_startofpacket     (alt_vip_cl_tpg_0_dout_startofpacket),                 //           .startofpacket
		.din_endofpacket       (alt_vip_cl_tpg_0_dout_endofpacket),                   //           .endofpacket
		.din_ready             (alt_vip_cl_tpg_0_dout_ready),                         //           .ready
		.dout_data             (main_scaler_dout_data),                               //       dout.data
		.dout_valid            (main_scaler_dout_valid),                              //           .valid
		.dout_startofpacket    (main_scaler_dout_startofpacket),                      //           .startofpacket
		.dout_endofpacket      (main_scaler_dout_endofpacket),                        //           .endofpacket
		.dout_ready            (main_scaler_dout_ready),                              //           .ready
		.control_address       (mm_interconnect_0_main_scaler_control_address),       //    control.address
		.control_byteenable    (mm_interconnect_0_main_scaler_control_byteenable),    //           .byteenable
		.control_write         (mm_interconnect_0_main_scaler_control_write),         //           .write
		.control_writedata     (mm_interconnect_0_main_scaler_control_writedata),     //           .writedata
		.control_read          (mm_interconnect_0_main_scaler_control_read),          //           .read
		.control_readdata      (mm_interconnect_0_main_scaler_control_readdata),      //           .readdata
		.control_readdatavalid (mm_interconnect_0_main_scaler_control_readdatavalid), //           .readdatavalid
		.control_waitrequest   (mm_interconnect_0_main_scaler_control_waitrequest)    //           .waitrequest
	);

	mySystem_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	mySystem_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	mySystem_pio_0 pio_0 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //                    .readdata
		.out_port   (pio_0_external_connection_export)       // external_connection.export
	);

	mySystem_uart_0 uart_0 (
		.clk           (clk_clk),                                   //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.rxd           (uart_0_external_connection_rxd),            // external_connection.export
		.txd           (uart_0_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver0_irq)                   //                 irq.irq
	);

	mySystem_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                    //                                clk_0_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                           //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                       //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                        //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                              //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                          //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                             //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                         //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                       //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                    //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                       //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                   //                                         .readdata
		.alt_vip_cl_mixer_0_control_address             (mm_interconnect_0_alt_vip_cl_mixer_0_control_address),       //               alt_vip_cl_mixer_0_control.address
		.alt_vip_cl_mixer_0_control_write               (mm_interconnect_0_alt_vip_cl_mixer_0_control_write),         //                                         .write
		.alt_vip_cl_mixer_0_control_read                (mm_interconnect_0_alt_vip_cl_mixer_0_control_read),          //                                         .read
		.alt_vip_cl_mixer_0_control_readdata            (mm_interconnect_0_alt_vip_cl_mixer_0_control_readdata),      //                                         .readdata
		.alt_vip_cl_mixer_0_control_writedata           (mm_interconnect_0_alt_vip_cl_mixer_0_control_writedata),     //                                         .writedata
		.alt_vip_cl_mixer_0_control_byteenable          (mm_interconnect_0_alt_vip_cl_mixer_0_control_byteenable),    //                                         .byteenable
		.alt_vip_cl_mixer_0_control_readdatavalid       (mm_interconnect_0_alt_vip_cl_mixer_0_control_readdatavalid), //                                         .readdatavalid
		.alt_vip_cl_mixer_0_control_waitrequest         (mm_interconnect_0_alt_vip_cl_mixer_0_control_waitrequest),   //                                         .waitrequest
		.alt_vip_cti_0_control_address                  (mm_interconnect_0_alt_vip_cti_0_control_address),            //                    alt_vip_cti_0_control.address
		.alt_vip_cti_0_control_write                    (mm_interconnect_0_alt_vip_cti_0_control_write),              //                                         .write
		.alt_vip_cti_0_control_read                     (mm_interconnect_0_alt_vip_cti_0_control_read),               //                                         .read
		.alt_vip_cti_0_control_readdata                 (mm_interconnect_0_alt_vip_cti_0_control_readdata),           //                                         .readdata
		.alt_vip_cti_0_control_writedata                (mm_interconnect_0_alt_vip_cti_0_control_writedata),          //                                         .writedata
		.main_scaler_control_address                    (mm_interconnect_0_main_scaler_control_address),              //                      main_scaler_control.address
		.main_scaler_control_write                      (mm_interconnect_0_main_scaler_control_write),                //                                         .write
		.main_scaler_control_read                       (mm_interconnect_0_main_scaler_control_read),                 //                                         .read
		.main_scaler_control_readdata                   (mm_interconnect_0_main_scaler_control_readdata),             //                                         .readdata
		.main_scaler_control_writedata                  (mm_interconnect_0_main_scaler_control_writedata),            //                                         .writedata
		.main_scaler_control_byteenable                 (mm_interconnect_0_main_scaler_control_byteenable),           //                                         .byteenable
		.main_scaler_control_readdatavalid              (mm_interconnect_0_main_scaler_control_readdatavalid),        //                                         .readdatavalid
		.main_scaler_control_waitrequest                (mm_interconnect_0_main_scaler_control_waitrequest),          //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),              //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),             //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),            //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),           //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),           //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                //                                         .clken
		.pio_0_s1_address                               (mm_interconnect_0_pio_0_s1_address),                         //                                 pio_0_s1.address
		.pio_0_s1_write                                 (mm_interconnect_0_pio_0_s1_write),                           //                                         .write
		.pio_0_s1_readdata                              (mm_interconnect_0_pio_0_s1_readdata),                        //                                         .readdata
		.pio_0_s1_writedata                             (mm_interconnect_0_pio_0_s1_writedata),                       //                                         .writedata
		.pio_0_s1_chipselect                            (mm_interconnect_0_pio_0_s1_chipselect),                      //                                         .chipselect
		.uart_0_s1_address                              (mm_interconnect_0_uart_0_s1_address),                        //                                uart_0_s1.address
		.uart_0_s1_write                                (mm_interconnect_0_uart_0_s1_write),                          //                                         .write
		.uart_0_s1_read                                 (mm_interconnect_0_uart_0_s1_read),                           //                                         .read
		.uart_0_s1_readdata                             (mm_interconnect_0_uart_0_s1_readdata),                       //                                         .readdata
		.uart_0_s1_writedata                            (mm_interconnect_0_uart_0_s1_writedata),                      //                                         .writedata
		.uart_0_s1_begintransfer                        (mm_interconnect_0_uart_0_s1_begintransfer),                  //                                         .begintransfer
		.uart_0_s1_chipselect                           (mm_interconnect_0_uart_0_s1_chipselect)                      //                                         .chipselect
	);

	mySystem_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                                                       (clk_clk),                                                                               //                                             clk_0_clk.clk
		.alt_vip_cl_vfb_0_mem_reset_reset_bridge_in_reset_reset              (rst_controller_reset_out_reset),                                                        //      alt_vip_cl_vfb_0_mem_reset_reset_bridge_in_reset.reset
		.alt_vip_cl_vfb_0_mem_master_rd_address                              (alt_vip_cl_vfb_0_mem_master_rd_address),                                                //                        alt_vip_cl_vfb_0_mem_master_rd.address
		.alt_vip_cl_vfb_0_mem_master_rd_waitrequest                          (alt_vip_cl_vfb_0_mem_master_rd_waitrequest),                                            //                                                      .waitrequest
		.alt_vip_cl_vfb_0_mem_master_rd_burstcount                           (alt_vip_cl_vfb_0_mem_master_rd_burstcount),                                             //                                                      .burstcount
		.alt_vip_cl_vfb_0_mem_master_rd_read                                 (alt_vip_cl_vfb_0_mem_master_rd_read),                                                   //                                                      .read
		.alt_vip_cl_vfb_0_mem_master_rd_readdata                             (alt_vip_cl_vfb_0_mem_master_rd_readdata),                                               //                                                      .readdata
		.alt_vip_cl_vfb_0_mem_master_rd_readdatavalid                        (alt_vip_cl_vfb_0_mem_master_rd_readdatavalid),                                          //                                                      .readdatavalid
		.alt_vip_cl_vfb_0_mem_master_wr_address                              (alt_vip_cl_vfb_0_mem_master_wr_address),                                                //                        alt_vip_cl_vfb_0_mem_master_wr.address
		.alt_vip_cl_vfb_0_mem_master_wr_waitrequest                          (alt_vip_cl_vfb_0_mem_master_wr_waitrequest),                                            //                                                      .waitrequest
		.alt_vip_cl_vfb_0_mem_master_wr_burstcount                           (alt_vip_cl_vfb_0_mem_master_wr_burstcount),                                             //                                                      .burstcount
		.alt_vip_cl_vfb_0_mem_master_wr_byteenable                           (alt_vip_cl_vfb_0_mem_master_wr_byteenable),                                             //                                                      .byteenable
		.alt_vip_cl_vfb_0_mem_master_wr_write                                (alt_vip_cl_vfb_0_mem_master_wr_write),                                                  //                                                      .write
		.alt_vip_cl_vfb_0_mem_master_wr_writedata                            (alt_vip_cl_vfb_0_mem_master_wr_writedata),                                              //                                                      .writedata
		.W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0_address       (mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_address),       // W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0.address
		.W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0_write         (mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_write),         //                                                      .write
		.W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0_read          (mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_read),          //                                                      .read
		.W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0_readdata      (mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_readdata),      //                                                      .readdata
		.W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0_writedata     (mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_writedata),     //                                                      .writedata
		.W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0_byteenable    (mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_byteenable),    //                                                      .byteenable
		.W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0_readdatavalid (mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_readdatavalid), //                                                      .readdatavalid
		.W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0_waitrequest   (mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_waitrequest),   //                                                      .waitrequest
		.W9825G6KH_SDRAMController_125MHz_CL3_0_avalon_slave_0_chipselect    (mm_interconnect_1_w9825g6kh_sdramcontroller_125mhz_cl3_0_avalon_slave_0_chipselect)     //                                                      .chipselect
	);

	mySystem_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
